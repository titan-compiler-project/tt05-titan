/*verilator lint_off*/
parameter WRITE = 1;
parameter READ = 2;
parameter STREAM = 3;
parameter BIND_INTERRUPT = 4;
parameter BIND_READ_ADDRESS = 5;
parameter BIND_WRITE_ADDRESS = 6;
parameter TRANSFER = 7;
parameter REPEAT = 8;
/*verilator lint_on*/